

module hoaaned_32b
(
  input [32-1:0] a,
  input [32-1:0] b,
  output [33-1:0] sum
);

  wire n1;
  wire n2;
  wire n3;
  wire n4;
  wire n5;
  wire cout12;
  wire cout16;
  wire cout20;
  wire cout24;
  wire cout28;
  assign sum[0] = 1;
  assign sum[1] = 1;
  assign sum[2] = 1;
  assign sum[3] = 1;
  assign sum[4] = 1;
  assign sum[5] = 1;
  assign sum[6] = 1;
  assign sum[7] = 1;

  or_2inp
  t1
  (
    .res(sum[8]),
    .inp1(a[8]),
    .inp2(b[8])
  );


  and_2inp
  t2
  (
    .res(n1),
    .inp1(a[8]),
    .inp2(b[8])
  );


  and_2inp
  t3
  (
    .res(n2),
    .inp1(a[9]),
    .inp2(b[9])
  );


  not_1inp
  t4
  (
    .res(n3),
    .inp(n2)
  );


  or_2inp
  t5
  (
    .res(n4),
    .inp1(a[9]),
    .inp2(b[9])
  );


  and_2inp
  t6
  (
    .res(n5),
    .inp1(n4),
    .inp2(n1)
  );


  or_2inp
  t7
  (
    .res(sum[9]),
    .inp1(n5),
    .inp2(n1)
  );


  frcla_2b
  cla1
  (
    .a1(a[11]),
    .a0(a[10]),
    .b1(b[11]),
    .b0(b[10]),
    .c0(n2),
    .c2(cout12),
    .sum1(sum[11]),
    .sum0(sum[10])
  );


  frcla_4b
  cla2
  (
    .a3(a[15]),
    .a2(a[14]),
    .a1(a[13]),
    .a0(a[12]),
    .b3(b[15]),
    .b2(b[14]),
    .b1(b[13]),
    .b0(b[12]),
    .c0(cout12),
    .c4(cout16),
    .sum3(sum[15]),
    .sum2(sum[14]),
    .sum1(sum[13]),
    .sum0(sum[12])
  );


  frcla_4b
  cla3
  (
    .a3(a[19]),
    .a2(a[18]),
    .a1(a[17]),
    .a0(a[16]),
    .b3(b[19]),
    .b2(b[18]),
    .b1(b[17]),
    .b0(b[16]),
    .c0(cout16),
    .c4(cout20),
    .sum3(sum[19]),
    .sum2(sum[18]),
    .sum1(sum[17]),
    .sum0(sum[16])
  );


  frcla_4b
  cla4
  (
    .a3(a[23]),
    .a2(a[22]),
    .a1(a[21]),
    .a0(a[20]),
    .b3(b[23]),
    .b2(b[22]),
    .b1(b[21]),
    .b0(b[20]),
    .c0(cout20),
    .c4(cout24),
    .sum3(sum[23]),
    .sum2(sum[22]),
    .sum1(sum[21]),
    .sum0(sum[20])
  );


  frcla_4b
  cla5
  (
    .a3(a[27]),
    .a2(a[26]),
    .a1(a[25]),
    .a0(a[24]),
    .b3(b[27]),
    .b2(b[26]),
    .b1(b[25]),
    .b0(b[24]),
    .c0(cout24),
    .c4(cout28),
    .sum3(sum[27]),
    .sum2(sum[26]),
    .sum1(sum[25]),
    .sum0(sum[24])
  );


  frcla_4b
  cla6
  (
    .a3(a[31]),
    .a2(a[30]),
    .a1(a[29]),
    .a0(a[28]),
    .b3(b[31]),
    .b2(b[30]),
    .b1(b[29]),
    .b0(b[28]),
    .c0(cout28),
    .c4(sum[32]),
    .sum3(sum[31]),
    .sum2(sum[30]),
    .sum1(sum[29]),
    .sum0(sum[28])
  );


endmodule



module or_2inp
(
  output res,
  input inp1,
  input inp2
);

  assign res = inp1 | inp2;

endmodule



module and_2inp
(
  output res,
  input inp1,
  input inp2
);

  assign res = inp1 & inp2;

endmodule



module not_1inp
(
  output res,
  input inp
);

  assign res = !inp;

endmodule



module frcla_2b
(
  input a1,
  input a0,
  input b1,
  input b0,
  input c0,
  output c2,
  output sum1,
  output sum0
);

  wire g1;
  wire g0;
  wire p1;
  wire p0;
  wire c1;
  wire m1;
  wire m2;

  and_2inp
  gate1
  (
    .res(g0),
    .inp1(a0),
    .inp2(b0)
  );


  and_2inp
  gate2
  (
    .res(g1),
    .inp1(a1),
    .inp2(b1)
  );


  xor_2inp
  gate5
  (
    .res(p0),
    .inp1(a0),
    .inp2(b0)
  );


  xor_2inp
  gate6
  (
    .res(p1),
    .inp1(a1),
    .inp2(b1)
  );


  ao21
  comp1
  (
    .a(p1),
    .b(g0),
    .c(g1),
    .y(m1)
  );


  and_2inp
  and1
  (
    .res(m2),
    .inp1(p1),
    .inp2(p0)
  );


  ao21
  comp6
  (
    .a(m2),
    .b(c0),
    .c(m1),
    .y(c2)
  );


  ao21
  comp7
  (
    .a(p0),
    .b(c0),
    .c(g0),
    .y(c1)
  );


  xor_2inp
  xorg1
  (
    .res(sum0),
    .inp1(p0),
    .inp2(c0)
  );


  xor_2inp
  xorg2
  (
    .res(sum1),
    .inp1(p1),
    .inp2(c1)
  );


endmodule



module xor_2inp
(
  output res,
  input inp1,
  input inp2
);

  assign res = inp1 ^ inp2;

endmodule



module ao21
(
  input a,
  input b,
  input c,
  output y
);

  wire net;

  and_2inp
  t1
  (
    .res(net),
    .inp1(a),
    .inp2(b)
  );


  or_2inp
  t2
  (
    .res(y),
    .inp1(net),
    .inp2(c)
  );


endmodule



module frcla_4b
(
  input a3,
  input a2,
  input a1,
  input a0,
  input b3,
  input b2,
  input b1,
  input b0,
  input c0,
  output c4,
  output sum3,
  output sum2,
  output sum1,
  output sum0
);

  wire g3;
  wire g2;
  wire g1;
  wire g0;
  wire p3;
  wire p2;
  wire p1;
  wire p0;
  wire c1;
  wire c2;
  wire c3;
  wire m1;
  wire m2;
  wire m3;
  wire m4;
  wire m5;
  wire m6;

  and_2inp
  gate1
  (
    .res(g0),
    .inp1(a0),
    .inp2(b0)
  );


  and_2inp
  gate2
  (
    .res(g1),
    .inp1(a1),
    .inp2(b1)
  );


  and_2inp
  gate3
  (
    .res(g2),
    .inp1(a2),
    .inp2(b2)
  );


  and_2inp
  gate4
  (
    .res(g3),
    .inp1(a3),
    .inp2(b3)
  );


  xor_2inp
  gate5
  (
    .res(p0),
    .inp1(a0),
    .inp2(b0)
  );


  xor_2inp
  gate6
  (
    .res(p1),
    .inp1(a1),
    .inp2(b1)
  );


  xor_2inp
  gate7
  (
    .res(p2),
    .inp1(a2),
    .inp2(b2)
  );


  xor_2inp
  gate8
  (
    .res(p3),
    .inp1(a3),
    .inp2(b3)
  );


  ao21
  comp1
  (
    .a(p1),
    .b(g0),
    .c(g1),
    .y(m1)
  );


  ao21
  comp2
  (
    .a(m1),
    .b(p2),
    .c(g2),
    .y(m2)
  );


  ao21
  comp3
  (
    .a(m2),
    .b(p3),
    .c(g3),
    .y(m3)
  );


  and_2inp
  and1
  (
    .res(m4),
    .inp1(p1),
    .inp2(p0)
  );


  and_2inp
  and2
  (
    .res(m5),
    .inp1(p2),
    .inp2(m4)
  );


  and_2inp
  and3
  (
    .res(m6),
    .inp1(p3),
    .inp2(m5)
  );


  ao21
  comp4
  (
    .a(m6),
    .b(c0),
    .c(m3),
    .y(c4)
  );


  ao21
  comp5
  (
    .a(m5),
    .b(c0),
    .c(m2),
    .y(c3)
  );


  ao21
  comp6
  (
    .a(m4),
    .b(c0),
    .c(m1),
    .y(c2)
  );


  ao21
  comp7
  (
    .a(p0),
    .b(c0),
    .c(g0),
    .y(c1)
  );


  xor_2inp
  xorg1
  (
    .res(sum0),
    .inp1(p0),
    .inp2(c0)
  );


  xor_2inp
  xorg2
  (
    .res(sum1),
    .inp1(p1),
    .inp2(c1)
  );


  xor_2inp
  xorg3
  (
    .res(sum2),
    .inp1(p2),
    .inp2(c2)
  );


  xor_2inp
  xorg4
  (
    .res(sum3),
    .inp1(p3),
    .inp2(c3)
  );


endmodule

